library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity MemoryM is
    Port(Data_In, Address : in STD_LOGIC_VECTOR(31 downto 0);
         MW : in STD_LOGIC;
         Data_Out : out STD_LOGIC_VECTOR(31 downto 0));
end MemoryM;

architecture Behavioral of MemoryM is
-- we will use the least significant 9 bit of the address - array(0 to 512)
type mem_array is array(0 to 511) of std_logic_vector(31 downto 0);
begin
mem_process: process (Address, Data_In)
variable data_mem : mem_array := (
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --  0 initialize processor i think
"00000000000" & "000001" & "00000" & "00000" & "00000", --  1 Fetch move mem
"00000000000" & "000001" & "00000" & "00000" & "00001", --  2 Fetch Move mem | Decode move 1 into reg0 
"00000000000" & "000011" & "00001" & "00000" & "00001", --  3 Fetch Add | Decode move 1 into reg1 | Execute move
"00000000000" & "000010" & "00000" & "00000" & "00001", --  4 Fetch move reg | decode add reg0 + reg1 -> reg0 | execute move
"00000000000" & "000100" & "00010" & "00000" & "00000", --  5 Fetch ADI | decode move reg 0 into reg2 | execute add
"00000000000" & "000101" & "00100" & "00000" & "00010", --  6 Fetch NOT | decode adI reg 0 + 2 -> reg4 | execute move
"00000000000" & "000110" & "00011" & "00000" & "00000", --  7 Fetch INC | decode not reg 0 -> reg3 | execute adi
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000111" & "00101" & "00000" & "00000", --  8 Fetch CMP | decode increment reg0 -> reg5 | execute not
"00000000000" & "001000" & "00000" & "00000" & "00000", --  9 Fetch BEQ | decode CMP reg0 and Reg 0 | execute INC
"00000000000" & "000011" & "00000" & "00000" & "00100", --  a Fetch B | decode offset to get to f = 4 | execute CMP
"00000000000" & "000011" & "00000" & "00000" & "00000", --  b Fetch ADD | Decode add reg 0+ reg0 -> reg0 | execute branch
"00000000000" & "000000" & "00000" & "00000" & "00000", --  c
"00000000000" & "000000" & "00000" & "00000" & "00000", --  d
"00000000000" & "000000" & "00000" & "00000" & "00000", --  e
"00000000000" & "001010" & "00000" & "00000" & "00000", --  f -Should branch here??? Fetch SR |
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "001011" & "00110" & "00000" & "00100", -- 10 Fetch B | deoce SR reg 4 -> reg 6
"00000000000" & "000001" & "00111" & "00000" & "01110", -- 11 Fetch X | decode branch offset -18 to 0 | execute SR
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 12 Fetch X | decode X | BRANCH
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 13 
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 14 
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 15
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 16
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 17
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 18
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 19
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 1a
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 1b
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 1c
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 1d
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 1e
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 1f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 20
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 21
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 22
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 23
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 24
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 25
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 26
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 27
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 28
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 29
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 2a
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 2b
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 2c
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 2d
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 2e
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 2f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 30
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 31
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 32
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 33
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 34
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 35
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 36
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 37
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 38
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 39
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 3a
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 3b
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 3c
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 3d
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 3e
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 3f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 40
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 41
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 42
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 43
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 44
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 45
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 46
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 47
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 48
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 49
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 4a
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 4b
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 4c
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 4d
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 4e
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 4f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 50
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 51
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 52
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 53
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 54
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 55
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 56
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 57
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 58
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 59
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 5a
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 5b
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 5c
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 5d
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 5e
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 5f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 60
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 61
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 62
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 63
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 64
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 65
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 66
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 67
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 68
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 69
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 6a
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 6b
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 6c
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 6d
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 6e
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 6f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 70
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 71
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 72
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 73
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 74
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 75
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 76
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 77
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 78
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 79
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 7a
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 7b
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 7c
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 7d
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 7e
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 7f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 80
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 81
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 82
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 83
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 84
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 85
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 86
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 87
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 88
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 89
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 8a
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 8b
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 8c
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 8d
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 8e
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 8f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 90
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 91
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 92
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 93
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 94
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 95
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 96
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 97
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 98
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 99
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 9a
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 9b
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 9c
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 9d
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 9e
"00000000000" & "000000" & "00000" & "00000" & "00000", -- 9f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- a0
"00000000000" & "000000" & "00000" & "00000" & "00000", -- a1
"00000000000" & "000000" & "00000" & "00000" & "00000", -- a2
"00000000000" & "000000" & "00000" & "00000" & "00000", -- a3
"00000000000" & "000000" & "00000" & "00000" & "00000", -- a4
"00000000000" & "000000" & "00000" & "00000" & "00000", -- a5
"00000000000" & "000000" & "00000" & "00000" & "00000", -- a6
"00000000000" & "000000" & "00000" & "00000" & "00000", -- a7
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- a8
"00000000000" & "000000" & "00000" & "00000" & "00000", -- a9
"00000000000" & "000000" & "00000" & "00000" & "00000", -- aa
"00000000000" & "000000" & "00000" & "00000" & "00000", -- ab
"00000000000" & "000000" & "00000" & "00000" & "00000", -- ac
"00000000000" & "000000" & "00000" & "00000" & "00000", -- ad
"00000000000" & "000000" & "00000" & "00000" & "00000", -- ae
"00000000000" & "000000" & "00000" & "00000" & "00000", -- af
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- b0
"00000000000" & "000000" & "00000" & "00000" & "00000", -- b1
"00000000000" & "000000" & "00000" & "00000" & "00000", -- b2
"00000000000" & "000000" & "00000" & "00000" & "00000", -- b3
"00000000000" & "000000" & "00000" & "00000" & "00000", -- b4
"00000000000" & "000000" & "00000" & "00000" & "00000", -- b5
"00000000000" & "000000" & "00000" & "00000" & "00000", -- b6
"00000000000" & "000000" & "00000" & "00000" & "00000", -- b7
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- b8
"00000000000" & "000000" & "00000" & "00000" & "00000", -- b9
"00000000000" & "000000" & "00000" & "00000" & "00000", -- ba
"00000000000" & "000000" & "00000" & "00000" & "00000", -- bb
"00000000000" & "000000" & "00000" & "00000" & "00000", -- bc
"00000000000" & "000000" & "00000" & "00000" & "00000", -- bd
"00000000000" & "000000" & "00000" & "00000" & "00000", -- be
"00000000000" & "000000" & "00000" & "00000" & "00000", -- bf
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- c0
"00000000000" & "000000" & "00000" & "00000" & "00000", -- c1
"00000000000" & "000000" & "00000" & "00000" & "00000", -- c2
"00000000000" & "000000" & "00000" & "00000" & "00000", -- c3
"00000000000" & "000000" & "00000" & "00000" & "00000", -- c4
"00000000000" & "000000" & "00000" & "00000" & "00000", -- c5
"00000000000" & "000000" & "00000" & "00000" & "00000", -- c6
"00000000000" & "000000" & "00000" & "00000" & "00000", -- c7
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- c8
"00000000000" & "000000" & "00000" & "00000" & "00000", -- c9
"00000000000" & "000000" & "00000" & "00000" & "00000", -- ca
"00000000000" & "000000" & "00000" & "00000" & "00000", -- cb
"00000000000" & "000000" & "00000" & "00000" & "00000", -- cc
"00000000000" & "000000" & "00000" & "00000" & "00000", -- cd
"00000000000" & "000000" & "00000" & "00000" & "00000", -- ce
"00000000000" & "000000" & "00000" & "00000" & "00000", -- cf
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- d0
"00000000000" & "000000" & "00000" & "00000" & "00000", -- d1
"00000000000" & "000000" & "00000" & "00000" & "00000", -- d2
"00000000000" & "000000" & "00000" & "00000" & "00000", -- d3
"00000000000" & "000000" & "00000" & "00000" & "00000", -- d4
"00000000000" & "000000" & "00000" & "00000" & "00000", -- d5
"00000000000" & "000000" & "00000" & "00000" & "00000", -- d6
"00000000000" & "000000" & "00000" & "00000" & "00000", -- d7
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- d8
"00000000000" & "000000" & "00000" & "00000" & "00000", -- d9
"00000000000" & "000000" & "00000" & "00000" & "00000", -- da
"00000000000" & "000000" & "00000" & "00000" & "00000", -- db
"00000000000" & "000000" & "00000" & "00000" & "00000", -- dc
"00000000000" & "000000" & "00000" & "00000" & "00000", -- dd
"00000000000" & "000000" & "00000" & "00000" & "00000", -- de
"00000000000" & "000000" & "00000" & "00000" & "00000", -- df
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- e0
"00000000000" & "000000" & "00000" & "00000" & "00000", -- e1
"00000000000" & "000000" & "00000" & "00000" & "00000", -- e2
"00000000000" & "000000" & "00000" & "00000" & "00000", -- e3
"00000000000" & "000000" & "00000" & "00000" & "00000", -- e4
"00000000000" & "000000" & "00000" & "00000" & "00000", -- e5
"00000000000" & "000000" & "00000" & "00000" & "00000", -- e6
"00000000000" & "000000" & "00000" & "00000" & "00000", -- e7
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- e8
"00000000000" & "000000" & "00000" & "00000" & "00000", -- e9
"00000000000" & "000000" & "00000" & "00000" & "00000", -- ea
"00000000000" & "000000" & "00000" & "00000" & "00000", -- eb
"00000000000" & "000000" & "00000" & "00000" & "00000", -- ec
"00000000000" & "000000" & "00000" & "00000" & "00000", -- ed
"00000000000" & "000000" & "00000" & "00000" & "00000", -- ee
"00000000000" & "000000" & "00000" & "00000" & "00000", -- ef
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- f0
"00000000000" & "000000" & "00000" & "00000" & "00000", -- f1
"00000000000" & "000000" & "00000" & "00000" & "00000", -- f2
"00000000000" & "000000" & "00000" & "00000" & "00000", -- f3
"00000000000" & "000000" & "00000" & "00000" & "00000", -- f4
"00000000000" & "000000" & "00000" & "00000" & "00000", -- f5
"00000000000" & "000000" & "00000" & "00000" & "00000", -- f6
"00000000000" & "000000" & "00000" & "00000" & "00000", -- f7
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", -- f8
"00000000000" & "000000" & "00000" & "00000" & "00000", -- f9
"00000000000" & "000000" & "00000" & "00000" & "00000", -- fa
"00000000000" & "000000" & "00000" & "00000" & "00000", -- fb
"00000000000" & "000000" & "00000" & "00000" & "00000", -- fc
"00000000000" & "000000" & "00000" & "00000" & "00000", -- fd
"00000000000" & "000000" & "00000" & "00000" & "00000", -- fe
"00000000000" & "000000" & "00000" & "00000" & "00000", -- ff
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --100
"00000000000" & "000000" & "00000" & "00000" & "00000", --101
"00000000000" & "000000" & "00000" & "00000" & "00000", --102
"00000000000" & "000000" & "00000" & "00000" & "00000", --103
"00000000000" & "000000" & "00000" & "00000" & "00000", --104
"00000000000" & "000000" & "00000" & "00000" & "00000", --105
"00000000000" & "000000" & "00000" & "00000" & "00000", --106
"00000000000" & "000000" & "00000" & "00000" & "00000", --107
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --108
"00000000000" & "000000" & "00000" & "00000" & "00000", --109
"00000000000" & "000000" & "00000" & "00000" & "00000", --10a
"00000000000" & "000000" & "00000" & "00000" & "00000", --10b
"00000000000" & "000000" & "00000" & "00000" & "00000", --10c
"00000000000" & "000000" & "00000" & "00000" & "00000", --10d
"00000000000" & "000000" & "00000" & "00000" & "00000", --10e
"00000000000" & "000000" & "00000" & "00000" & "00000", --10f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --110
"00000000000" & "000000" & "00000" & "00000" & "00000", --111
"00000000000" & "000000" & "00000" & "00000" & "00000", --112
"00000000000" & "000000" & "00000" & "00000" & "00000", --113
"00000000000" & "000000" & "00000" & "00000" & "00000", --114
"00000000000" & "000000" & "00000" & "00000" & "00000", --115
"00000000000" & "000000" & "00000" & "00000" & "00000", --116
"00000000000" & "000000" & "00000" & "00000" & "00000", --117
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --118
"00000000000" & "000000" & "00000" & "00000" & "00000", --119
"00000000000" & "000000" & "00000" & "00000" & "00000", --11a
"00000000000" & "000000" & "00000" & "00000" & "00000", --11b
"00000000000" & "000000" & "00000" & "00000" & "00000", --11c
"00000000000" & "000000" & "00000" & "00000" & "00000", --11d
"00000000000" & "000000" & "00000" & "00000" & "00000", --11e
"00000000000" & "000000" & "00000" & "00000" & "00000", --11f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --120
"00000000000" & "000000" & "00000" & "00000" & "00000", --121
"00000000000" & "000000" & "00000" & "00000" & "00000", --122
"00000000000" & "000000" & "00000" & "00000" & "00000", --123
"00000000000" & "000000" & "00000" & "00000" & "00000", --124
"00000000000" & "000000" & "00000" & "00000" & "00000", --125
"00000000000" & "000000" & "00000" & "00000" & "00000", --126
"00000000000" & "000000" & "00000" & "00000" & "00000", --127
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --128
"00000000000" & "000000" & "00000" & "00000" & "00000", --129
"00000000000" & "000000" & "00000" & "00000" & "00000", --12a
"00000000000" & "000000" & "00000" & "00000" & "00000", --12b
"00000000000" & "000000" & "00000" & "00000" & "00000", --12c
"00000000000" & "000000" & "00000" & "00000" & "00000", --12d
"00000000000" & "000000" & "00000" & "00000" & "00000", --12e
"00000000000" & "000000" & "00000" & "00000" & "00000", --12f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --130
"00000000000" & "000000" & "00000" & "00000" & "00000", --131
"00000000000" & "000000" & "00000" & "00000" & "00000", --132
"00000000000" & "000000" & "00000" & "00000" & "00000", --133
"00000000000" & "000000" & "00000" & "00000" & "00000", --134
"00000000000" & "000000" & "00000" & "00000" & "00000", --135
"00000000000" & "000000" & "00000" & "00000" & "00000", --136
"00000000000" & "000000" & "00000" & "00000" & "00000", --137
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --138
"00000000000" & "000000" & "00000" & "00000" & "00000", --139
"00000000000" & "000000" & "00000" & "00000" & "00000", --13a
"00000000000" & "000000" & "00000" & "00000" & "00000", --13b
"00000000000" & "000000" & "00000" & "00000" & "00000", --13c
"00000000000" & "000000" & "00000" & "00000" & "00000", --13d
"00000000000" & "000000" & "00000" & "00000" & "00000", --13e
"00000000000" & "000000" & "00000" & "00000" & "00000", --13f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --140
"00000000000" & "000000" & "00000" & "00000" & "00000", --141
"00000000000" & "000000" & "00000" & "00000" & "00000", --142
"00000000000" & "000000" & "00000" & "00000" & "00000", --143
"00000000000" & "000000" & "00000" & "00000" & "00000", --144
"00000000000" & "000000" & "00000" & "00000" & "00000", --145
"00000000000" & "000000" & "00000" & "00000" & "00000", --146
"00000000000" & "000000" & "00000" & "00000" & "00000", --147
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --148
"00000000000" & "000000" & "00000" & "00000" & "00000", --149
"00000000000" & "000000" & "00000" & "00000" & "00000", --14a
"00000000000" & "000000" & "00000" & "00000" & "00000", --14b
"00000000000" & "000000" & "00000" & "00000" & "00000", --14c
"00000000000" & "000000" & "00000" & "00000" & "00000", --14d
"00000000000" & "000000" & "00000" & "00000" & "00000", --14e
"00000000000" & "000000" & "00000" & "00000" & "00000", --14f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --150
"00000000000" & "000000" & "00000" & "00000" & "00000", --151
"00000000000" & "000000" & "00000" & "00000" & "00000", --152
"00000000000" & "000000" & "00000" & "00000" & "00000", --153
"00000000000" & "000000" & "00000" & "00000" & "00000", --154
"00000000000" & "000000" & "00000" & "00000" & "00000", --155
"00000000000" & "000000" & "00000" & "00000" & "00000", --156
"00000000000" & "000000" & "00000" & "00000" & "00000", --157
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --158
"00000000000" & "000000" & "00000" & "00000" & "00000", --159
"00000000000" & "000000" & "00000" & "00000" & "00000", --15a
"00000000000" & "000000" & "00000" & "00000" & "00000", --15b
"00000000000" & "000000" & "00000" & "00000" & "00000", --15c
"00000000000" & "000000" & "00000" & "00000" & "00000", --15d
"00000000000" & "000000" & "00000" & "00000" & "00000", --15e
"00000000000" & "000000" & "00000" & "00000" & "00000", --15f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --160
"00000000000" & "000000" & "00000" & "00000" & "00000", --161
"00000000000" & "000000" & "00000" & "00000" & "00000", --162
"00000000000" & "000000" & "00000" & "00000" & "00000", --163
"00000000000" & "000000" & "00000" & "00000" & "00000", --164
"00000000000" & "000000" & "00000" & "00000" & "00000", --165
"00000000000" & "000000" & "00000" & "00000" & "00000", --166
"00000000000" & "000000" & "00000" & "00000" & "00000", --167
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --168
"00000000000" & "000000" & "00000" & "00000" & "00000", --169
"00000000000" & "000000" & "00000" & "00000" & "00000", --16a
"00000000000" & "000000" & "00000" & "00000" & "00000", --16b
"00000000000" & "000000" & "00000" & "00000" & "00000", --16c
"00000000000" & "000000" & "00000" & "00000" & "00000", --16d
"00000000000" & "000000" & "00000" & "00000" & "00000", --16e
"00000000000" & "000000" & "00000" & "00000" & "00000", --16f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --170
"00000000000" & "000000" & "00000" & "00000" & "00000", --171
"00000000000" & "000000" & "00000" & "00000" & "00000", --172
"00000000000" & "000000" & "00000" & "00000" & "00000", --173
"00000000000" & "000000" & "00000" & "00000" & "00000", --174
"00000000000" & "000000" & "00000" & "00000" & "00000", --175
"00000000000" & "000000" & "00000" & "00000" & "00000", --176
"00000000000" & "000000" & "00000" & "00000" & "00000", --177
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --178
"00000000000" & "000000" & "00000" & "00000" & "00000", --179
"00000000000" & "000000" & "00000" & "00000" & "00000", --17a
"00000000000" & "000000" & "00000" & "00000" & "00000", --17b
"00000000000" & "000000" & "00000" & "00000" & "00000", --17c
"00000000000" & "000000" & "00000" & "00000" & "00000", --17d
"00000000000" & "000000" & "00000" & "00000" & "00000", --17e
"00000000000" & "000000" & "00000" & "00000" & "00000", --17f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --180
"00000000000" & "000000" & "00000" & "00000" & "00000", --181
"00000000000" & "000000" & "00000" & "00000" & "00000", --182
"00000000000" & "000000" & "00000" & "00000" & "00000", --183
"00000000000" & "000000" & "00000" & "00000" & "00000", --184
"00000000000" & "000000" & "00000" & "00000" & "00000", --185
"00000000000" & "000000" & "00000" & "00000" & "00000", --186
"00000000000" & "000000" & "00000" & "00000" & "00000", --187
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --188
"00000000000" & "000000" & "00000" & "00000" & "00000", --189
"00000000000" & "000000" & "00000" & "00000" & "00000", --18a
"00000000000" & "000000" & "00000" & "00000" & "00000", --18b
"00000000000" & "000000" & "00000" & "00000" & "00000", --18c
"00000000000" & "000000" & "00000" & "00000" & "00000", --18d
"00000000000" & "000000" & "00000" & "00000" & "00000", --18e
"00000000000" & "000000" & "00000" & "00000" & "00000", --18f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --190
"00000000000" & "000000" & "00000" & "00000" & "00000", --191
"00000000000" & "000000" & "00000" & "00000" & "00000", --192
"00000000000" & "000000" & "00000" & "00000" & "00000", --193
"00000000000" & "000000" & "00000" & "00000" & "00000", --194
"00000000000" & "000000" & "00000" & "00000" & "00000", --195
"00000000000" & "000000" & "00000" & "00000" & "00000", --196
"00000000000" & "000000" & "00000" & "00000" & "00000", --197
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --198
"00000000000" & "000000" & "00000" & "00000" & "00000", --199
"00000000000" & "000000" & "00000" & "00000" & "00000", --19a
"00000000000" & "000000" & "00000" & "00000" & "00000", --19b
"00000000000" & "000000" & "00000" & "00000" & "00000", --19c
"00000000000" & "000000" & "00000" & "00000" & "00000", --19d
"00000000000" & "000000" & "00000" & "00000" & "00000", --19e
"00000000000" & "000000" & "00000" & "00000" & "00000", --19f
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --1a0
"00000000000" & "000000" & "00000" & "00000" & "00000", --1a1
"00000000000" & "000000" & "00000" & "00000" & "00000", --1a2
"00000000000" & "000000" & "00000" & "00000" & "00000", --1a3
"00000000000" & "000000" & "00000" & "00000" & "00000", --1a4
"00000000000" & "000000" & "00000" & "00000" & "00000", --1a5
"00000000000" & "000000" & "00000" & "00000" & "00000", --1a6
"00000000000" & "000000" & "00000" & "00000" & "00000", --1a7
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --1a8
"00000000000" & "000000" & "00000" & "00000" & "00000", --1a9
"00000000000" & "000000" & "00000" & "00000" & "00000", --1aa
"00000000000" & "000000" & "00000" & "00000" & "00000", --1ab
"00000000000" & "000000" & "00000" & "00000" & "00000", --1ac
"00000000000" & "000000" & "00000" & "00000" & "00000", --1ad
"00000000000" & "000000" & "00000" & "00000" & "00000", --1ae
"00000000000" & "000000" & "00000" & "00000" & "00000", --1af
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --1b0
"00000000000" & "000000" & "00000" & "00000" & "00000", --1b1
"00000000000" & "000000" & "00000" & "00000" & "00000", --1b2
"00000000000" & "000000" & "00000" & "00000" & "00000", --1b3
"00000000000" & "000000" & "00000" & "00000" & "00000", --1b4
"00000000000" & "000000" & "00000" & "00000" & "00000", --1b5
"00000000000" & "000000" & "00000" & "00000" & "00000", --1b6
"00000000000" & "000000" & "00000" & "00000" & "00000", --1b7
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --1b8
"00000000000" & "000000" & "00000" & "00000" & "00000", --1b9
"00000000000" & "000000" & "00000" & "00000" & "00000", --1ba
"00000000000" & "000000" & "00000" & "00000" & "00000", --1bb
"00000000000" & "000000" & "00000" & "00000" & "00000", --1bc
"00000000000" & "000000" & "00000" & "00000" & "00000", --1bd
"00000000000" & "000000" & "00000" & "00000" & "00000", --1be
"00000000000" & "000000" & "00000" & "00000" & "00000", --1bf
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --1c0
"00000000000" & "000000" & "00000" & "00000" & "00000", --1c1
"00000000000" & "000000" & "00000" & "00000" & "00000", --1c2
"00000000000" & "000000" & "00000" & "00000" & "00000", --1c3
"00000000000" & "000000" & "00000" & "00000" & "00000", --1c4
"00000000000" & "000000" & "00000" & "00000" & "00000", --1c5
"00000000000" & "000000" & "00000" & "00000" & "00000", --1c6
"00000000000" & "000000" & "00000" & "00000" & "00000", --1c7
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --1c8
"00000000000" & "000000" & "00000" & "00000" & "00000", --1c9
"00000000000" & "000000" & "00000" & "00000" & "00000", --1ca
"00000000000" & "000000" & "00000" & "00000" & "00000", --1cb
"00000000000" & "000000" & "00000" & "00000" & "00000", --1cc
"00000000000" & "000000" & "00000" & "00000" & "00000", --1cd
"00000000000" & "000000" & "00000" & "00000" & "00000", --1ce
"00000000000" & "000000" & "00000" & "00000" & "00000", --1cf
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --1d0
"00000000000" & "000000" & "00000" & "00000" & "00000", --1d1
"00000000000" & "000000" & "00000" & "00000" & "00000", --1d2
"00000000000" & "000000" & "00000" & "00000" & "00000", --1d3
"00000000000" & "000000" & "00000" & "00000" & "00000", --1d4
"00000000000" & "000000" & "00000" & "00000" & "00000", --1d5
"00000000000" & "000000" & "00000" & "00000" & "00000", --1d6
"00000000000" & "000000" & "00000" & "00000" & "00000", --1d7
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --1d8
"00000000000" & "000000" & "00000" & "00000" & "00000", --1d9
"00000000000" & "000000" & "00000" & "00000" & "00000", --1da
"00000000000" & "000000" & "00000" & "00000" & "00000", --1db
"00000000000" & "000000" & "00000" & "00000" & "00000", --1dc
"00000000000" & "000000" & "00000" & "00000" & "00000", --1dd
"00000000000" & "000000" & "00000" & "00000" & "00000", --1de
"00000000000" & "000000" & "00000" & "00000" & "00000", --1df
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --1e0
"00000000000" & "000000" & "00000" & "00000" & "00000", --1e1
"00000000000" & "000000" & "00000" & "00000" & "00000", --1e2
"00000000000" & "000000" & "00000" & "00000" & "00000", --1e3
"00000000000" & "000000" & "00000" & "00000" & "00000", --1e4
"00000000000" & "000000" & "00000" & "00000" & "00000", --1e5
"00000000000" & "000000" & "00000" & "00000" & "00000", --1e6
"00000000000" & "000000" & "00000" & "00000" & "00000", --1e7
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --1e8
"00000000000" & "000000" & "00000" & "00000" & "00000", --1e9
"00000000000" & "000000" & "00000" & "00000" & "00000", --1ea
"00000000000" & "000000" & "00000" & "00000" & "00000", --1eb
"00000000000" & "000000" & "00000" & "00000" & "00000", --1ec
"00000000000" & "000000" & "00000" & "00000" & "00000", --1ed
"00000000000" & "000000" & "00000" & "00000" & "00000", --1ee
"00000000000" & "000000" & "00000" & "00000" & "00000", --1ef
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --1f0
"00000000000" & "000000" & "00000" & "00000" & "00000", --1f1
"00000000000" & "000000" & "00000" & "00000" & "00000", --1f2
"00000000000" & "000000" & "00000" & "00000" & "00000", --1f3
"00000000000" & "000000" & "00000" & "00000" & "00000", --1f4
"00000000000" & "000000" & "00000" & "00000" & "00000", --1f5
"00000000000" & "000000" & "00000" & "00000" & "00000", --1f6
"00000000000" & "000000" & "00000" & "00000" & "00000", --1f7
--| Not Used |  OpCode  |    DR   |    SA   |   SB   |
"00000000000" & "000000" & "00000" & "00000" & "00000", --1f8
"00000000000" & "000000" & "00000" & "00000" & "00000", --1f9
"00000000000" & "000000" & "00000" & "00000" & "00000", --1fa
"00000000000" & "000000" & "00000" & "00000" & "00000", --1fb
"00000000000" & "000000" & "00000" & "00000" & "00000", --1fc
"00000000000" & "000000" & "00000" & "00000" & "00000", --1fd
"00000000000" & "000000" & "00000" & "00000" & "00000", --1fe
"00000000000" & "000000" & "00000" & "00000" & "00000" --1ff
);
variable addr : integer;
begin -- the following type conversion function is in std_logic_arith
addr := conv_integer(unsigned(Address(8 downto 0)));

if MW ='1' then
data_mem(addr):= Data_In;
end if;
Data_Out <= data_mem(addr) after 10 ns;

end process;
end Behavioral;


