library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity OldDecoder5To32 is
    Port ( 
     DestA : in std_logic_vector(4 downto 0);
     DestChoice : out std_logic_vector(31 downto 0));    
end OldDecoder5To32;

architecture Behavioral of OldDecoder5To32 is
begin
with DestA select
DestChoice <= "00000000000000000000000000000001" after 5ns when "00000",
              "00000000000000000000000000000010" after 5ns when "00001",
              "00000000000000000000000000000100" after 5ns when "00010",
              "00000000000000000000000000001000" after 5ns when "00011",
              "00000000000000000000000000010000" after 5ns when "00100",
              "00000000000000000000000000100000" after 5ns when "00101",
              "00000000000000000000000001000000" after 5ns when "00110",
              "00000000000000000000000010000000" after 5ns when "00111",
              "00000000000000000000000100000000" after 5ns when "01000",
              "00000000000000000000001000000000" after 5ns when "01001",
              "00000000000000000000010000000000" after 5ns when "01010",
              "00000000000000000000100000000000" after 5ns when "01011",
              "00000000000000000001000000000000" after 5ns when "01100",
              "00000000000000000010000000000000" after 5ns when "01101",
              "00000000000000000100000000000000" after 5ns when "01110",
              "00000000000000001000000000000000" after 5ns when "01111",
              "00000000000000010000000000000000" after 5ns when "10000",
              "00000000000000100000000000000000" after 5ns when "10001",
              "00000000000001000000000000000000" after 5ns when "10010",
              "00000000000010000000000000000000" after 5ns when "10011",
              "00000000000100000000000000000000" after 5ns when "10100",
              "00000000001000000000000000000000" after 5ns when "10101",
              "00000000010000000000000000000000" after 5ns when "10110",
              "00000000100000000000000000000000" after 5ns when "10111",
              "00000001000000000000000000000000" after 5ns when "11000",
              "00000010000000000000000000000000" after 5ns when "11001",
              "00000100000000000000000000000000" after 5ns when "11010",
              "00001000000000000000000000000000" after 5ns when "11011",
              "00010000000000000000000000000000" after 5ns when "11100",
              "00100000000000000000000000000000" after 5ns when "11101",
              "01000000000000000000000000000000" after 5ns when "11110",
              "10000000000000000000000000000000" after 5ns when "11111",
              "00000000000000000000000000000000" when others;
end Behavioral;
