library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MUX32_5_32TB is
end MUX32_5_32TB;

architecture Behavioral of MUX32_5_32TB is
    component MUX32_5_32 
        Port(
          R00, R01, R02, R03, R04, R05, R06, R07, R08, R09 ,R10, R11, R12, R13, R14, R15, R16, R17, R18, R19, R20, R21, R22 ,R23, R24, R25, R26, R27, R28, R29, R30, R31, R32 : in STD_LOGIC_VECTOR(31 downto 0);
          S : in STD_LOGIC_VECTOR (4 downto 0);
          T : in STD_LOGIC;
          DataOut : out STD_LOGIC_VECTOR (31 downto 0));
    end component;
    
    signal R00, R01, R02, R03, R04, R05 : STD_LOGIC_VECTOR(31 downto 0);
    signal R06, R07, R08, R09 ,R10, R11 : STD_LOGIC_VECTOR(31 downto 0);
    signal R12, R13, R14, R15, R16, R17 : STD_LOGIC_VECTOR(31 downto 0);
    signal R18, R19, R20, R21, R22 ,R23 : STD_LOGIC_VECTOR(31 downto 0);
    signal R24, R25, R26, R27, R28, R29 : STD_LOGIC_VECTOR(31 downto 0);
    signal R30, R31, R32 : STD_LOGIC_VECTOR(31 downto 0);
    signal T : STD_LOGIC;
    signal S : STD_LOGIC_VECTOR (4 downto 0);
    signal DataOut : STD_LOGIC_VECTOR (31 downto 0);
begin
UUT : MUX32_5_32 port map(R00 => R00, R01 => R01, R02 => R02, R03 => R03, R04 => R04, R05 => R05, R06 => R06, R07 => R07, R08 => R08, R09 => R09,R10 => R10, R11 => R11, R12 => R12, R13 => R13, R14 => R14, R15 => R15, R16 => R16, R17 => R17, R18 => R18, R19 => R19,R20 => R20, R21 => R21, R22 => R22, R23 => R23, R24 => R24, R25 => R25, R26 => R26, R27 => R27, R28 => R28, R29 => R29,R30 => R30, R31 => R31, R32 => R32, S => S,  T => T, DataOut => DataOut);
Multi3232_run : process
    begin
        R00 <= "00000000000000000000000000000001";
        R01 <= "00000000000000000000000000000010";
        R02 <= "00000000000000000000000000000100";
        R03 <= "00000000000000000000000000001000";
        R04 <= "00000000000000000000000000010000";
        R05 <= "00000000000000000000000000100000";
        R06 <= "00000000000000000000000001000000";
        R07 <= "00000000000000000000000010000000";
        R08 <= "00000000000000000000000100000000";
        R09 <= "00000000000000000000001000000000";
        R10 <= "00000000000000000000010000000000";
        R11 <= "00000000000000000000100000000000";
        R12 <= "00000000000000000001000000000000";
        R13 <= "00000000000000000010000000000000";
        R14 <= "00000000000000000100000000000000";
        R15 <= "00000000000000001000000000000000";
        R16 <= "00000000000000010000000000000000";
        R17 <= "00000000000000100000000000000000";
        R18 <= "00000000000001000000000000000000";
        R19 <= "00000000000010000000000000000000";
        R20 <= "00000000000100000000000000000000";
        R21 <= "00000000001000000000000000000000";
        R22 <= "00000000010000000000000000000000";
        R23 <= "00000000100000000000000000000000";
        R24 <= "00000001000000000000000000000000";
        R25 <= "00000010000000000000000000000000";
        R26 <= "00000100000000000000000000000000";
        R27 <= "00001000000000000000000000000000";
        R28 <= "00010000000000000000000000000000";
        R29 <= "00100000000000000000000000000000";
        R30 <= "01000000000000000000000000000000";
        R31 <= "10000000000000000000000000000000";
        R32 <= "11111111111111111111111111111111";
        
        T <= '0';
        S <= "00000";
        wait for 10ns;
        S <= "00001";
        wait for 10ns;
        S <= "00010";
        wait for 10ns;
        S <= "00011";
        wait for 10ns;
        S <= "00100";
        wait for 10ns;
        S <= "00101";
        wait for 10ns;
        S <= "00110";
        wait for 10ns;
        S <= "00111";
        wait for 10ns;
        S <= "01000";
        wait for 10ns;
        S <= "01001";
        wait for 10ns;
        S <= "01010";
        wait for 10ns;
        S <= "01011";
        wait for 10ns;
        S <= "01100";
        wait for 10ns;
        S <= "01101";
        wait for 10ns;
        S <= "01110";
        wait for 10ns;
        S <= "01111";
        wait for 10ns;
        S <= "10000";
        wait for 10ns;
        S <= "10001";
        wait for 10ns;
        S <= "10010";
        wait for 10ns;
        S <= "10011";
        wait for 10ns;
        S <= "10100";
        wait for 10ns;
        S <= "10101";
        wait for 10ns;
        S <= "10110";
        wait for 10ns;
        S <= "10111";
        wait for 10ns;
        S <= "11000";
        wait for 10ns;
        S <= "11001";
        wait for 10ns;
        S <= "11010";
        wait for 10ns;
        S <= "11011";
        wait for 10ns;
        S <= "11100";
        wait for 10ns;
        S <= "11101";
        wait for 10ns;
        S <= "11110";
        wait for 10ns;
        S <= "11111";
        wait for 10ns;
        T <= '1';
        wait for 10ns;
      
     end process;       
end Behavioral;
